
module Video_change (
	probe,
	source_clk,
	source);	

	input	[31:0]	probe;
	input		source_clk;
	output	[31:0]	source;
endmodule

// cram_clock_en.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module cram_clock_en (
		input  wire  inclk,  //  altclkctrl_input.inclk
		input  wire  ena,    //                  .ena
		output wire  outclk  // altclkctrl_output.outclk
	);

	cram_clock_en_altclkctrl_0 altclkctrl_0 (
		.inclk  (inclk),  //  altclkctrl_input.inclk
		.ena    (ena),    //                  .ena
		.outclk (outclk)  // altclkctrl_output.outclk
	);

endmodule

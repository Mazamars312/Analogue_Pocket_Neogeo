//
// microrom and nanorom instantiation
//
// There is bit of wasting of resources here. An extra registering pipeline happens that is not needed.
// This is just for the purpose of helping inferring block RAM using pure generic code. Inferring RAM is important for performance.
// Might be more efficient to use vendor specific features such as clock enable.
//

module uRom( input clk, input [UADDR_WIDTH-1:0] microAddr, output reg [UROM_WIDTH-1:0] microOutput);
	reg [UROM_WIDTH-1:0] uRam[ UROM_DEPTH];		
	initial begin
uRam[0   ] <= 17'b10010000101100000;
uRam[1   ] <= 17'b10000100000000000;
uRam[2   ] <= 17'b00101001011010000;
uRam[3   ] <= 17'b00111110011000000;
uRam[4   ] <= 17'b01000000000001100;
uRam[5   ] <= 17'b01000000000001100;
uRam[6   ] <= 17'b01000010010000000;
uRam[7   ] <= 17'b10001100011100000;
uRam[8   ] <= 17'b01000100010000000;
uRam[9   ] <= 17'b10000000010000000;
uRam[10  ] <= 17'b10000000010000000;
uRam[11  ] <= 17'b01000100010000000;
uRam[12  ] <= 17'b00001010010000000;
uRam[13  ] <= 17'b10000000100000000;
uRam[14  ] <= 17'b10000000100000000;
uRam[15  ] <= 17'b01101001100000000;
uRam[16  ] <= 17'b00000000000000000;
uRam[17  ] <= 17'b00000000000000000;
uRam[18  ] <= 17'b00000000000000000;
uRam[19  ] <= 17'b00000000000000000;
uRam[20  ] <= 17'b00000000000000000;
uRam[21  ] <= 17'b00000000000000000;
uRam[22  ] <= 17'b00000000000000000;
uRam[23  ] <= 17'b00000000000000000;
uRam[24  ] <= 17'b00000000000000000;
uRam[25  ] <= 17'b00000000000000000;
uRam[26  ] <= 17'b00000000000000000;
uRam[27  ] <= 17'b00000000000000000;
uRam[28  ] <= 17'b00000000000000000;
uRam[29  ] <= 17'b00000000000000000;
uRam[30  ] <= 17'b00000000000000000;
uRam[31  ] <= 17'b00000000000000000;
uRam[32  ] <= 17'b00000000000000100;
uRam[33  ] <= 17'b00001010110000000;
uRam[34  ] <= 17'b00111000001100000;
uRam[35  ] <= 17'b00100101001001010;
uRam[36  ] <= 17'b00000000000001100;
uRam[37  ] <= 17'b10110000110100001;
uRam[38  ] <= 17'b00000000000001100;
uRam[39  ] <= 17'b00001110100000000;
uRam[40  ] <= 17'b00110100101000000;
uRam[41  ] <= 17'b00100011010100000;
uRam[42  ] <= 17'b00000010010000000;
uRam[43  ] <= 17'b10000110000000010;
uRam[44  ] <= 17'b00111110110000000;
uRam[45  ] <= 17'b00000100011100000;
uRam[46  ] <= 17'b00101111010100000;
uRam[47  ] <= 17'b10010011100000010;
uRam[48  ] <= 17'b00000000000000000;
uRam[49  ] <= 17'b00000000000000000;
uRam[50  ] <= 17'b00000000000000000;
uRam[51  ] <= 17'b00000000000000000;
uRam[52  ] <= 17'b00000000000000000;
uRam[53  ] <= 17'b00000000000000000;
uRam[54  ] <= 17'b00000000000000000;
uRam[55  ] <= 17'b00000000000000000;
uRam[56  ] <= 17'b00000000000000000;
uRam[57  ] <= 17'b00000000000000000;
uRam[58  ] <= 17'b00000000000000000;
uRam[59  ] <= 17'b00000000000000000;
uRam[60  ] <= 17'b00000000000000000;
uRam[61  ] <= 17'b00000000000000000;
uRam[62  ] <= 17'b00000000000000000;
uRam[63  ] <= 17'b00000000000000000;
uRam[64  ] <= 17'b10011101000000000;
uRam[65  ] <= 17'b00000100110010110;
uRam[66  ] <= 17'b00101001010000000;
uRam[67  ] <= 17'b10110000110100001;
uRam[68  ] <= 17'b00000000000000100;
uRam[69  ] <= 17'b00111110000100000;
uRam[70  ] <= 17'b10010111010100000;
uRam[71  ] <= 17'b01000110000100000;
uRam[72  ] <= 17'b01010111100000000;
uRam[73  ] <= 17'b10001010010011010;
uRam[74  ] <= 17'b01000110010100001;
uRam[75  ] <= 17'b00000110010111010;
uRam[76  ] <= 17'b01001100010100000;
uRam[77  ] <= 17'b10001010010010111;
uRam[78  ] <= 17'b01000000000100001;
uRam[79  ] <= 17'b00110100111000000;
uRam[80  ] <= 17'b00000000000000000;
uRam[81  ] <= 17'b00000000000000000;
uRam[82  ] <= 17'b00000000000000000;
uRam[83  ] <= 17'b00000000000000000;
uRam[84  ] <= 17'b00000000000000000;
uRam[85  ] <= 17'b00000000000000000;
uRam[86  ] <= 17'b00000000000000000;
uRam[87  ] <= 17'b00000000000000000;
uRam[88  ] <= 17'b00000000000000000;
uRam[89  ] <= 17'b00000000000000000;
uRam[90  ] <= 17'b00000000000000000;
uRam[91  ] <= 17'b00000000000000000;
uRam[92  ] <= 17'b00000000000000000;
uRam[93  ] <= 17'b00000000000000000;
uRam[94  ] <= 17'b00000000000000000;
uRam[95  ] <= 17'b00000000000000000;
uRam[96  ] <= 17'b00000010001100000;
uRam[97  ] <= 17'b01001010000100001;
uRam[98  ] <= 17'b10110100111000000;
uRam[99  ] <= 17'b00011011010100000;
uRam[100 ] <= 17'b10000000000000100;
uRam[101 ] <= 17'b10110100111000000;
uRam[102 ] <= 17'b00000000000000100;
uRam[103 ] <= 17'b00001000001000000;
uRam[104 ] <= 17'b00000100011100110;
uRam[105 ] <= 17'b10001110010100001;
uRam[106 ] <= 17'b00000000011110010;
uRam[107 ] <= 17'b01001000011000000;
uRam[108 ] <= 17'b00001000010100110;
uRam[109 ] <= 17'b10001010000110111;
uRam[110 ] <= 17'b00000000111110010;
uRam[111 ] <= 17'b01001000111000000;
uRam[112 ] <= 17'b00000000000000000;
uRam[113 ] <= 17'b00000000000000000;
uRam[114 ] <= 17'b00000000000000000;
uRam[115 ] <= 17'b00000000000000000;
uRam[116 ] <= 17'b00000000000000000;
uRam[117 ] <= 17'b00000000000000000;
uRam[118 ] <= 17'b00000000000000000;
uRam[119 ] <= 17'b00000000000000000;
uRam[120 ] <= 17'b00000000000000000;
uRam[121 ] <= 17'b00000000000000000;
uRam[122 ] <= 17'b00000000000000000;
uRam[123 ] <= 17'b00000000000000000;
uRam[124 ] <= 17'b00000000000000000;
uRam[125 ] <= 17'b00000000000000000;
uRam[126 ] <= 17'b00000000000000000;
uRam[127 ] <= 17'b00000000000000000;
uRam[128 ] <= 17'b10101001000000001;
uRam[129 ] <= 17'b10001000001000001;
uRam[130 ] <= 17'b01000000000000100;
uRam[131 ] <= 17'b01001100001111010;
uRam[132 ] <= 17'b00000110001000000;
uRam[133 ] <= 17'b00010110001100000;
uRam[134 ] <= 17'b00011010000000000;
uRam[135 ] <= 17'b10110000110100001;
uRam[136 ] <= 17'b01111000001100000;
uRam[137 ] <= 17'b00011000000000000;
uRam[138 ] <= 17'b00000100100100001;
uRam[139 ] <= 17'b00000000000000100;
uRam[140 ] <= 17'b00000000101100000;
uRam[141 ] <= 17'b00000000000000100;
uRam[142 ] <= 17'b00010001010100000;
uRam[143 ] <= 17'b10010111000100001;
uRam[144 ] <= 17'b00000000000000000;
uRam[145 ] <= 17'b00000000000000000;
uRam[146 ] <= 17'b00000000000000000;
uRam[147 ] <= 17'b00000000000000000;
uRam[148 ] <= 17'b00000000000000000;
uRam[149 ] <= 17'b00000000000000000;
uRam[150 ] <= 17'b00000000000000000;
uRam[151 ] <= 17'b00000000000000000;
uRam[152 ] <= 17'b00000000000000000;
uRam[153 ] <= 17'b00000000000000000;
uRam[154 ] <= 17'b00000000000000000;
uRam[155 ] <= 17'b00000000000000000;
uRam[156 ] <= 17'b00000000000000000;
uRam[157 ] <= 17'b00000000000000000;
uRam[158 ] <= 17'b00000000000000000;
uRam[159 ] <= 17'b00000000000000000;
uRam[160 ] <= 17'b00000010001100000;
uRam[161 ] <= 17'b00000000000000100;
uRam[162 ] <= 17'b01111000011100000;
uRam[163 ] <= 17'b00011011010100000;
uRam[164 ] <= 17'b00101101000000000;
uRam[165 ] <= 17'b01000110010111010;
uRam[166 ] <= 17'b00101101000000000;
uRam[167 ] <= 17'b10001010101100000;
uRam[168 ] <= 17'b01010110001100000;
uRam[169 ] <= 17'b00011000110000000;
uRam[170 ] <= 17'b01010110001100000;
uRam[171 ] <= 17'b10001110011100001;
uRam[172 ] <= 17'b00000100101100000;
uRam[173 ] <= 17'b01000110010111010;
uRam[174 ] <= 17'b00000100101100000;
uRam[175 ] <= 17'b10001010111100000;
uRam[176 ] <= 17'b00000000000000000;
uRam[177 ] <= 17'b00000000000000000;
uRam[178 ] <= 17'b00000000000000000;
uRam[179 ] <= 17'b00000000000000000;
uRam[180 ] <= 17'b00000000000000000;
uRam[181 ] <= 17'b00000000000000000;
uRam[182 ] <= 17'b00000000000000000;
uRam[183 ] <= 17'b00000000000000000;
uRam[184 ] <= 17'b00000000000000000;
uRam[185 ] <= 17'b00000000000000000;
uRam[186 ] <= 17'b00000000000000000;
uRam[187 ] <= 17'b00000000000000000;
uRam[188 ] <= 17'b00000000000000000;
uRam[189 ] <= 17'b00000000000000000;
uRam[190 ] <= 17'b00000000000000000;
uRam[191 ] <= 17'b00000000000000000;
uRam[192 ] <= 17'b10101001000000001;
uRam[193 ] <= 17'b00001000101010110;
uRam[194 ] <= 17'b00011111010100000;
uRam[195 ] <= 17'b01101101110000000;
uRam[196 ] <= 17'b00000000000000100;
uRam[197 ] <= 17'b10111110000100000;
uRam[198 ] <= 17'b00000100011100000;
uRam[199 ] <= 17'b10001100101000001;
uRam[200 ] <= 17'b00000110001000000;
uRam[201 ] <= 17'b00001110000010010;
uRam[202 ] <= 17'b00100101000010110;
uRam[203 ] <= 17'b00101101000100000;
uRam[204 ] <= 17'b00000000011100000;
uRam[205 ] <= 17'b00001000111100000;
uRam[206 ] <= 17'b00100101000011010;
uRam[207 ] <= 17'b00110100111000000;
uRam[208 ] <= 17'b00000000000000000;
uRam[209 ] <= 17'b00000000000000000;
uRam[210 ] <= 17'b00000000000000000;
uRam[211 ] <= 17'b00000000000000000;
uRam[212 ] <= 17'b00000000000000000;
uRam[213 ] <= 17'b00000000000000000;
uRam[214 ] <= 17'b00000000000000000;
uRam[215 ] <= 17'b00000000000000000;
uRam[216 ] <= 17'b00000000000000000;
uRam[217 ] <= 17'b00000000000000000;
uRam[218 ] <= 17'b00000000000000000;
uRam[219 ] <= 17'b00000000000000000;
uRam[220 ] <= 17'b00000000000000000;
uRam[221 ] <= 17'b00000000000000000;
uRam[222 ] <= 17'b00000000000000000;
uRam[223 ] <= 17'b00000000000000000;
uRam[224 ] <= 17'b00000010000100010;
uRam[225 ] <= 17'b00001010110000000;
uRam[226 ] <= 17'b00000000000000100;
uRam[227 ] <= 17'b00101101010000000;
uRam[228 ] <= 17'b01010001010000000;
uRam[229 ] <= 17'b01000110111000000;
uRam[230 ] <= 17'b00000000000000100;
uRam[231 ] <= 17'b00000000010110010;
uRam[232 ] <= 17'b00110100101000000;
uRam[233 ] <= 17'b00100011010100000;
uRam[234 ] <= 17'b10000000000001000;
uRam[235 ] <= 17'b01101011010000000;
uRam[236 ] <= 17'b00111110110000000;
uRam[237 ] <= 17'b00000100011100000;
uRam[238 ] <= 17'b10010101000000000;
uRam[239 ] <= 17'b01111110010100000;
uRam[240 ] <= 17'b00000000000000000;
uRam[241 ] <= 17'b00000000000000000;
uRam[242 ] <= 17'b00000000000000000;
uRam[243 ] <= 17'b00000000000000000;
uRam[244 ] <= 17'b00000000000000000;
uRam[245 ] <= 17'b00000000000000000;
uRam[246 ] <= 17'b00000000000000000;
uRam[247 ] <= 17'b00000000000000000;
uRam[248 ] <= 17'b00000000000000000;
uRam[249 ] <= 17'b00000000000000000;
uRam[250 ] <= 17'b00000000000000000;
uRam[251 ] <= 17'b00000000000000000;
uRam[252 ] <= 17'b00000000000000000;
uRam[253 ] <= 17'b00000000000000000;
uRam[254 ] <= 17'b00000000000000000;
uRam[255 ] <= 17'b00000000000000000;
uRam[256 ] <= 17'b10001100101000001;
uRam[257 ] <= 17'b10000010100000010;
uRam[258 ] <= 17'b01000010101000000;
uRam[259 ] <= 17'b00011111100100000;
uRam[260 ] <= 17'b10100111100000001;
uRam[261 ] <= 17'b10010010110000010;
uRam[262 ] <= 17'b01110100111000000;
uRam[263 ] <= 17'b00010111010000000;
uRam[264 ] <= 17'b10101011100000001;
uRam[265 ] <= 17'b10010010100000010;
uRam[266 ] <= 17'b01110000100100000;
uRam[267 ] <= 17'b00000000100100000;
uRam[268 ] <= 17'b10100101100100001;
uRam[269 ] <= 17'b10000010110000010;
uRam[270 ] <= 17'b01001010101000000;
uRam[271 ] <= 17'b00010111000000000;
uRam[272 ] <= 17'b00010001000010110;
uRam[273 ] <= 17'b01110010100111010;
uRam[274 ] <= 17'b10110100010000000;
uRam[275 ] <= 17'b00110100111000000;
uRam[276 ] <= 17'b01000010010000110;
uRam[277 ] <= 17'b01110010110111011;
uRam[278 ] <= 17'b01111100000000000;
uRam[279 ] <= 17'b00101101000100000;
uRam[280 ] <= 17'b00101001001010001;
uRam[281 ] <= 17'b01011011111100000;
uRam[282 ] <= 17'b01101111011000000;
uRam[283 ] <= 17'b00100011100000000;
uRam[284 ] <= 17'b00111110000110000;
uRam[285 ] <= 17'b00000000000000000;
uRam[286 ] <= 17'b10101111011000000;
uRam[287 ] <= 17'b00000000000000000;
uRam[288 ] <= 17'b00001010100000000;
uRam[289 ] <= 17'b10101011100100001;
uRam[290 ] <= 17'b01010011000100001;
uRam[291 ] <= 17'b10010101010000000;
uRam[292 ] <= 17'b00000000110000000;
uRam[293 ] <= 17'b10111010000100001;
uRam[294 ] <= 17'b01011001010000000;
uRam[295 ] <= 17'b10010101000000000;
uRam[296 ] <= 17'b00101101101100000;
uRam[297 ] <= 17'b10100011100100001;
uRam[298 ] <= 17'b01011110100000000;
uRam[299 ] <= 17'b01110100011100000;
uRam[300 ] <= 17'b00101011111000000;
uRam[301 ] <= 17'b10110000110100001;
uRam[302 ] <= 17'b01010101010100001;
uRam[303 ] <= 17'b00000000000000000;
uRam[304 ] <= 17'b00111000100000000;
uRam[305 ] <= 17'b01011011000000000;
uRam[306 ] <= 17'b00001000100100000;
uRam[307 ] <= 17'b10001100101000001;
uRam[308 ] <= 17'b00100001100000000;
uRam[309 ] <= 17'b01011011010000000;
uRam[310 ] <= 17'b00001000110100000;
uRam[311 ] <= 17'b10011001110100001;
uRam[312 ] <= 17'b00000110010111010;
uRam[313 ] <= 17'b01011011100000000;
uRam[314 ] <= 17'b00000000110100000;
uRam[315 ] <= 17'b10011101010000001;
uRam[316 ] <= 17'b00000000000000000;
uRam[317 ] <= 17'b00000000000000000;
uRam[318 ] <= 17'b00000000000000000;
uRam[319 ] <= 17'b00000000000000000;
uRam[320 ] <= 17'b00000000000000000;
uRam[321 ] <= 17'b00000000000000000;
uRam[322 ] <= 17'b00000000000000000;
uRam[323 ] <= 17'b00000000000000000;
uRam[324 ] <= 17'b00000000000000000;
uRam[325 ] <= 17'b00000000000000000;
uRam[326 ] <= 17'b00000000000000000;
uRam[327 ] <= 17'b00000000000000000;
uRam[328 ] <= 17'b00000000000000000;
uRam[329 ] <= 17'b00000000000000000;
uRam[330 ] <= 17'b00000000000000000;
uRam[331 ] <= 17'b00000000000000000;
uRam[332 ] <= 17'b00000000000000000;
uRam[333 ] <= 17'b00000000000000000;
uRam[334 ] <= 17'b00000000000000000;
uRam[335 ] <= 17'b00000000000000000;
uRam[336 ] <= 17'b10110000110100001;
uRam[337 ] <= 17'b00011101000100000;
uRam[338 ] <= 17'b00011101000100000;
uRam[339 ] <= 17'b00010001000101110;
uRam[340 ] <= 17'b01011010110000000;
uRam[341 ] <= 17'b01011001010100000;
uRam[342 ] <= 17'b10011101010100000;
uRam[343 ] <= 17'b00000000000000100;
uRam[344 ] <= 17'b10110000110100001;
uRam[345 ] <= 17'b00110110000000000;
uRam[346 ] <= 17'b10110000011100001;
uRam[347 ] <= 17'b10110000011100001;
uRam[348 ] <= 17'b10011101000000001;
uRam[349 ] <= 17'b01110100111000000;
uRam[350 ] <= 17'b00101101100100000;
uRam[351 ] <= 17'b10011000100000000;
uRam[352 ] <= 17'b00000000000000000;
uRam[353 ] <= 17'b00000000000000000;
uRam[354 ] <= 17'b00000000000000000;
uRam[355 ] <= 17'b00000000000000000;
uRam[356 ] <= 17'b00000000000000000;
uRam[357 ] <= 17'b00000000000000000;
uRam[358 ] <= 17'b00000000000000000;
uRam[359 ] <= 17'b00000000000000000;
uRam[360 ] <= 17'b00000000000000000;
uRam[361 ] <= 17'b00000000000000000;
uRam[362 ] <= 17'b00000000000000000;
uRam[363 ] <= 17'b00000000000000000;
uRam[364 ] <= 17'b00000000000000000;
uRam[365 ] <= 17'b00000000000000000;
uRam[366 ] <= 17'b00000000000000000;
uRam[367 ] <= 17'b00000000000000000;
uRam[368 ] <= 17'b10000000000000100;
uRam[369 ] <= 17'b00000000000000100;
uRam[370 ] <= 17'b00000100111000000;
uRam[371 ] <= 17'b00000100111000000;
uRam[372 ] <= 17'b00000100111000000;
uRam[373 ] <= 17'b00001100010101010;
uRam[374 ] <= 17'b00001000000010110;
uRam[375 ] <= 17'b00101001010000000;
uRam[376 ] <= 17'b10011000100000000;
uRam[377 ] <= 17'b00011011100100000;
uRam[378 ] <= 17'b01000100010000000;
uRam[379 ] <= 17'b01000000000001100;
uRam[380 ] <= 17'b10011000010000001;
uRam[381 ] <= 17'b10011011110100000;
uRam[382 ] <= 17'b10011111110100001;
uRam[383 ] <= 17'b00011000010000000;
uRam[384 ] <= 17'b00000000000000000;
uRam[385 ] <= 17'b00000000000000000;
uRam[386 ] <= 17'b00000000000000000;
uRam[387 ] <= 17'b00000000000000000;
uRam[388 ] <= 17'b00000000000000000;
uRam[389 ] <= 17'b00000000000000000;
uRam[390 ] <= 17'b00000000000000000;
uRam[391 ] <= 17'b00000000000000000;
uRam[392 ] <= 17'b00000000000000000;
uRam[393 ] <= 17'b00000000000000000;
uRam[394 ] <= 17'b00000000000000000;
uRam[395 ] <= 17'b00000000000000000;
uRam[396 ] <= 17'b00000000000000000;
uRam[397 ] <= 17'b00000000000000000;
uRam[398 ] <= 17'b00000000000000000;
uRam[399 ] <= 17'b00000000000000000;
uRam[400 ] <= 17'b00000000000000000;
uRam[401 ] <= 17'b00000000000000000;
uRam[402 ] <= 17'b00000000000000000;
uRam[403 ] <= 17'b00000000000000000;
uRam[404 ] <= 17'b00000000000000000;
uRam[405 ] <= 17'b00000000000000000;
uRam[406 ] <= 17'b00000000000000000;
uRam[407 ] <= 17'b00000000000000000;
uRam[408 ] <= 17'b00000000000000000;
uRam[409 ] <= 17'b00000000000000000;
uRam[410 ] <= 17'b00000000000000000;
uRam[411 ] <= 17'b00000000000000000;
uRam[412 ] <= 17'b00000000000000000;
uRam[413 ] <= 17'b00000000000000000;
uRam[414 ] <= 17'b00000000000000000;
uRam[415 ] <= 17'b00000000000000000;
uRam[416 ] <= 17'b00000000000000000;
uRam[417 ] <= 17'b00000000000000000;
uRam[418 ] <= 17'b00000000000000000;
uRam[419 ] <= 17'b00000000000000000;
uRam[420 ] <= 17'b00000000000000000;
uRam[421 ] <= 17'b00000000000000000;
uRam[422 ] <= 17'b00000000000000000;
uRam[423 ] <= 17'b00000000000000000;
uRam[424 ] <= 17'b00000000000000000;
uRam[425 ] <= 17'b00000000000000000;
uRam[426 ] <= 17'b00000000000000000;
uRam[427 ] <= 17'b00000000000000000;
uRam[428 ] <= 17'b00000000000000000;
uRam[429 ] <= 17'b00000000000000000;
uRam[430 ] <= 17'b00000000000000000;
uRam[431 ] <= 17'b00000000000000000;
uRam[432 ] <= 17'b00000000000000000;
uRam[433 ] <= 17'b00000000000000000;
uRam[434 ] <= 17'b00000000000000000;
uRam[435 ] <= 17'b00000000000000000;
uRam[436 ] <= 17'b00000000000000000;
uRam[437 ] <= 17'b00000000000000000;
uRam[438 ] <= 17'b00000000000000000;
uRam[439 ] <= 17'b00000000000000000;
uRam[440 ] <= 17'b00000000000000000;
uRam[441 ] <= 17'b00000000000000000;
uRam[442 ] <= 17'b00000000000000000;
uRam[443 ] <= 17'b00000000000000000;
uRam[444 ] <= 17'b00000000000000000;
uRam[445 ] <= 17'b00000000000000000;
uRam[446 ] <= 17'b00000000000000000;
uRam[447 ] <= 17'b00000000000000000;
uRam[448 ] <= 17'b00111110001000000;
uRam[449 ] <= 17'b10101011100100001;
uRam[450 ] <= 17'b10001010100000000;
uRam[451 ] <= 17'b10101011100100001;
uRam[452 ] <= 17'b00100011010000000;
uRam[453 ] <= 17'b10110000001100001;
uRam[454 ] <= 17'b10000000110000000;
uRam[455 ] <= 17'b10110000101100001;
uRam[456 ] <= 17'b00000000000000000;
uRam[457 ] <= 17'b10110000101100001;
uRam[458 ] <= 17'b10110110110100000;
uRam[459 ] <= 17'b10100001110100001;
uRam[460 ] <= 17'b00111100010000000;
uRam[461 ] <= 17'b10011101100000001;
uRam[462 ] <= 17'b10111110100100000;
uRam[463 ] <= 17'b10010011010100001;
uRam[464 ] <= 17'b00111100010100000;
uRam[465 ] <= 17'b10101011100000001;
uRam[466 ] <= 17'b10101001101000000;
uRam[467 ] <= 17'b10101011100000001;
uRam[468 ] <= 17'b00000000000000000;
uRam[469 ] <= 17'b10011111000100001;
uRam[470 ] <= 17'b10101001111000000;
uRam[471 ] <= 17'b10011011000100001;
uRam[472 ] <= 17'b00000000000000000;
uRam[473 ] <= 17'b10010011010100001;
uRam[474 ] <= 17'b00000000000000000;
uRam[475 ] <= 17'b00000000000000000;
uRam[476 ] <= 17'b00000000000000000;
uRam[477 ] <= 17'b00000000000000000;
uRam[478 ] <= 17'b00000000000000000;
uRam[479 ] <= 17'b00000000000000000;
uRam[480 ] <= 17'b00001010100000000;
uRam[481 ] <= 17'b10111110000100000;
uRam[482 ] <= 17'b10000100100000000;
uRam[483 ] <= 17'b00111010001100000;
uRam[484 ] <= 17'b00000000110000000;
uRam[485 ] <= 17'b10011001000000000;
uRam[486 ] <= 17'b10000100110000000;
uRam[487 ] <= 17'b00111010011100000;
uRam[488 ] <= 17'b00101101101100000;
uRam[489 ] <= 17'b10001110111000000;
uRam[490 ] <= 17'b10101111101000000;
uRam[491 ] <= 17'b00010100100000000;
uRam[492 ] <= 17'b00101011111000000;
uRam[493 ] <= 17'b10110100001100000;
uRam[494 ] <= 17'b10101111111000000;
uRam[495 ] <= 17'b00010100010000000;
uRam[496 ] <= 17'b00111000100000000;
uRam[497 ] <= 17'b10110100101100000;
uRam[498 ] <= 17'b10101001010100000;
uRam[499 ] <= 17'b00101011001000000;
uRam[500 ] <= 17'b00100001100000000;
uRam[501 ] <= 17'b10001110010000000;
uRam[502 ] <= 17'b10101111001000000;
uRam[503 ] <= 17'b00101011011000000;
uRam[504 ] <= 17'b00000110010111010;
uRam[505 ] <= 17'b10111000110000000;
uRam[506 ] <= 17'b10011101110100000;
uRam[507 ] <= 17'b00111010101100000;
uRam[508 ] <= 17'b00000000000000000;
uRam[509 ] <= 17'b10101011011100000;
uRam[510 ] <= 17'b01100011110100001;
uRam[511 ] <= 17'b00111010111100000;
uRam[512 ] <= 17'b00000000000000000;
uRam[513 ] <= 17'b00000000000000000;
uRam[514 ] <= 17'b00000000000000000;
uRam[515 ] <= 17'b00000000000000000;
uRam[516 ] <= 17'b00000000000000000;
uRam[517 ] <= 17'b00000000000000000;
uRam[518 ] <= 17'b00000000000000000;
uRam[519 ] <= 17'b00000000000000000;
uRam[520 ] <= 17'b00000000000000000;
uRam[521 ] <= 17'b00000000000000000;
uRam[522 ] <= 17'b00000000000000000;
uRam[523 ] <= 17'b00000000000000000;
uRam[524 ] <= 17'b00000000000000000;
uRam[525 ] <= 17'b00000000000000000;
uRam[526 ] <= 17'b00000000000000000;
uRam[527 ] <= 17'b00000000000000000;
uRam[528 ] <= 17'b00100101000000000;
uRam[529 ] <= 17'b00000100000010110;
uRam[530 ] <= 17'b00000000000000100;
uRam[531 ] <= 17'b00001110000001110;
uRam[532 ] <= 17'b00100001000000000;
uRam[533 ] <= 17'b10110000110100001;
uRam[534 ] <= 17'b00100101011001010;
uRam[535 ] <= 17'b00111000001100000;
uRam[536 ] <= 17'b00100101100000001;
uRam[537 ] <= 17'b10011000010000000;
uRam[538 ] <= 17'b01101101100000000;
uRam[539 ] <= 17'b00000000000001100;
uRam[540 ] <= 17'b01100101110000000;
uRam[541 ] <= 17'b00000000000001100;
uRam[542 ] <= 17'b00001100001111010;
uRam[543 ] <= 17'b01001100001111010;
uRam[544 ] <= 17'b00000000000000000;
uRam[545 ] <= 17'b00000000000000000;
uRam[546 ] <= 17'b00000000000000000;
uRam[547 ] <= 17'b00000000000000000;
uRam[548 ] <= 17'b00000000000000000;
uRam[549 ] <= 17'b00000000000000000;
uRam[550 ] <= 17'b00000000000000000;
uRam[551 ] <= 17'b00000000000000000;
uRam[552 ] <= 17'b00000000000000000;
uRam[553 ] <= 17'b00000000000000000;
uRam[554 ] <= 17'b00000000000000000;
uRam[555 ] <= 17'b00000000000000000;
uRam[556 ] <= 17'b00000000000000000;
uRam[557 ] <= 17'b00000000000000000;
uRam[558 ] <= 17'b00000000000000000;
uRam[559 ] <= 17'b00000000000000000;
uRam[560 ] <= 17'b10101111000000001;
uRam[561 ] <= 17'b00000100111000000;
uRam[562 ] <= 17'b10101111000000001;
uRam[563 ] <= 17'b00000000000000100;
uRam[564 ] <= 17'b00100111010000000;
uRam[565 ] <= 17'b00001110101100000;
uRam[566 ] <= 17'b11010001100000000;
uRam[567 ] <= 17'b00110010100111010;
uRam[568 ] <= 17'b00000000000000100;
uRam[569 ] <= 17'b00000100111000000;
uRam[570 ] <= 17'b00000000000000100;
uRam[571 ] <= 17'b10110000110100001;
uRam[572 ] <= 17'b01100111110000001;
uRam[573 ] <= 17'b10000000000000100;
uRam[574 ] <= 17'b01111100100100000;
uRam[575 ] <= 17'b01100001100100001;
uRam[576 ] <= 17'b00000000000000000;
uRam[577 ] <= 17'b00000000000000000;
uRam[578 ] <= 17'b00000000000000000;
uRam[579 ] <= 17'b00000000000000000;
uRam[580 ] <= 17'b00000000000000000;
uRam[581 ] <= 17'b00000000000000000;
uRam[582 ] <= 17'b00000000000000000;
uRam[583 ] <= 17'b00000000000000000;
uRam[584 ] <= 17'b00000000000000000;
uRam[585 ] <= 17'b00000000000000000;
uRam[586 ] <= 17'b00000000000000000;
uRam[587 ] <= 17'b00000000000000000;
uRam[588 ] <= 17'b00000000000000000;
uRam[589 ] <= 17'b00000000000000000;
uRam[590 ] <= 17'b00000000000000000;
uRam[591 ] <= 17'b00000000000000000;
uRam[592 ] <= 17'b00000000001100000;
uRam[593 ] <= 17'b10001010010100001;
uRam[594 ] <= 17'b00110110100000110;
uRam[595 ] <= 17'b00000000000000100;
uRam[596 ] <= 17'b00100001000000000;
uRam[597 ] <= 17'b10111110000100000;
uRam[598 ] <= 17'b10100111000100000;
uRam[599 ] <= 17'b00111000010000000;
uRam[600 ] <= 17'b10000000000000100;
uRam[601 ] <= 17'b00101001100100000;
uRam[602 ] <= 17'b00101101100100000;
uRam[603 ] <= 17'b00000000000000100;
uRam[604 ] <= 17'b00100101110100000;
uRam[605 ] <= 17'b00000000000000100;
uRam[606 ] <= 17'b00100101110100000;
uRam[607 ] <= 17'b00100101110100000;
uRam[608 ] <= 17'b00000000000000000;
uRam[609 ] <= 17'b00000000000000000;
uRam[610 ] <= 17'b00000000000000000;
uRam[611 ] <= 17'b00000000000000000;
uRam[612 ] <= 17'b00000000000000000;
uRam[613 ] <= 17'b00000000000000000;
uRam[614 ] <= 17'b00000000000000000;
uRam[615 ] <= 17'b00000000000000000;
uRam[616 ] <= 17'b00000000000000000;
uRam[617 ] <= 17'b00000000000000000;
uRam[618 ] <= 17'b00000000000000000;
uRam[619 ] <= 17'b00000000000000000;
uRam[620 ] <= 17'b00000000000000000;
uRam[621 ] <= 17'b00000000000000000;
uRam[622 ] <= 17'b00000000000000000;
uRam[623 ] <= 17'b00000000000000000;
uRam[624 ] <= 17'b10100111000100000;
uRam[625 ] <= 17'b01101011000100000;
uRam[626 ] <= 17'b01111110000100001;
uRam[627 ] <= 17'b10100111000100000;
uRam[628 ] <= 17'b10100111001000000;
uRam[629 ] <= 17'b10111110000100000;
uRam[630 ] <= 17'b00101111010000000;
uRam[631 ] <= 17'b00110010100111010;
uRam[632 ] <= 17'b00000000000000100;
uRam[633 ] <= 17'b10100011100100001;
uRam[634 ] <= 17'b00000000000000100;
uRam[635 ] <= 17'b00000010011100001;
uRam[636 ] <= 17'b10100111110100000;
uRam[637 ] <= 17'b00000000000000100;
uRam[638 ] <= 17'b00101111110100000;
uRam[639 ] <= 17'b00101111101100000;
uRam[640 ] <= 17'b00000000000000000;
uRam[641 ] <= 17'b00000000000000000;
uRam[642 ] <= 17'b00000000000000000;
uRam[643 ] <= 17'b00000000000000000;
uRam[644 ] <= 17'b00000000000000000;
uRam[645 ] <= 17'b00000000000000000;
uRam[646 ] <= 17'b00000000000000000;
uRam[647 ] <= 17'b00000000000000000;
uRam[648 ] <= 17'b00000000000000000;
uRam[649 ] <= 17'b00000000000000000;
uRam[650 ] <= 17'b00000000000000000;
uRam[651 ] <= 17'b00000000000000000;
uRam[652 ] <= 17'b00000000000000000;
uRam[653 ] <= 17'b00000000000000000;
uRam[654 ] <= 17'b00000000000000000;
uRam[655 ] <= 17'b00000000000000000;
uRam[656 ] <= 17'b00100101001000000;
uRam[657 ] <= 17'b00101001000010110;
uRam[658 ] <= 17'b00110010000100000;
uRam[659 ] <= 17'b00100011000100000;
uRam[660 ] <= 17'b00100101011000000;
uRam[661 ] <= 17'b00101001011100000;
uRam[662 ] <= 17'b00101011110110000;
uRam[663 ] <= 17'b00101111001000000;
uRam[664 ] <= 17'b00010100000000000;
uRam[665 ] <= 17'b10110100111000001;
uRam[666 ] <= 17'b01110010100100000;
uRam[667 ] <= 17'b10110000110100001;
uRam[668 ] <= 17'b00010100110000000;
uRam[669 ] <= 17'b10110100110100001;
uRam[670 ] <= 17'b01111000110100000;
uRam[671 ] <= 17'b10111110110100001;
uRam[672 ] <= 17'b00000000000000000;
uRam[673 ] <= 17'b00000000000000000;
uRam[674 ] <= 17'b00000000000000000;
uRam[675 ] <= 17'b00000000000000000;
uRam[676 ] <= 17'b00000000000000000;
uRam[677 ] <= 17'b00000000000000000;
uRam[678 ] <= 17'b00000000000000000;
uRam[679 ] <= 17'b00000000000000000;
uRam[680 ] <= 17'b00000000000000000;
uRam[681 ] <= 17'b00000000000000000;
uRam[682 ] <= 17'b00000000000000000;
uRam[683 ] <= 17'b00000000000000000;
uRam[684 ] <= 17'b00000000000000000;
uRam[685 ] <= 17'b00000000000000000;
uRam[686 ] <= 17'b00000000000000000;
uRam[687 ] <= 17'b00000000000000000;
uRam[688 ] <= 17'b00100011010100000;
uRam[689 ] <= 17'b00100111000100000;
uRam[690 ] <= 17'b00000110100000010;
uRam[691 ] <= 17'b10111110000100000;
uRam[692 ] <= 17'b00000100011100000;
uRam[693 ] <= 17'b00110000110000000;
uRam[694 ] <= 17'b00000110110000010;
uRam[695 ] <= 17'b10010001110000000;
uRam[696 ] <= 17'b10110100111000001;
uRam[697 ] <= 17'b10000000000001000;
uRam[698 ] <= 17'b01110000100100000;
uRam[699 ] <= 17'b10110100101000000;
uRam[700 ] <= 17'b10010101110100001;
uRam[701 ] <= 17'b10111110000100000;
uRam[702 ] <= 17'b01101101111100000;
uRam[703 ] <= 17'b10101011101000000;
uRam[704 ] <= 17'b00000000000000000;
uRam[705 ] <= 17'b00000000000000000;
uRam[706 ] <= 17'b00000000000000000;
uRam[707 ] <= 17'b00000000000000000;
uRam[708 ] <= 17'b00000000000000000;
uRam[709 ] <= 17'b00000000000000000;
uRam[710 ] <= 17'b00000000000000000;
uRam[711 ] <= 17'b00000000000000000;
uRam[712 ] <= 17'b00000000000000000;
uRam[713 ] <= 17'b00000000000000000;
uRam[714 ] <= 17'b00000000000000000;
uRam[715 ] <= 17'b00000000000000000;
uRam[716 ] <= 17'b00000000000000000;
uRam[717 ] <= 17'b00000000000000000;
uRam[718 ] <= 17'b00000000000000000;
uRam[719 ] <= 17'b00000000000000000;
uRam[720 ] <= 17'b00101001000010110;
uRam[721 ] <= 17'b10001010011100001;
uRam[722 ] <= 17'b00100001000000110;
uRam[723 ] <= 17'b00101101000000110;
uRam[724 ] <= 17'b00101001011100000;
uRam[725 ] <= 17'b10001010011100001;
uRam[726 ] <= 17'b00110110111000110;
uRam[727 ] <= 17'b00101101010000110;
uRam[728 ] <= 17'b10001100101000001;
uRam[729 ] <= 17'b10110100101000000;
uRam[730 ] <= 17'b10101101101100000;
uRam[731 ] <= 17'b01111110000100001;
uRam[732 ] <= 17'b10100101100100001;
uRam[733 ] <= 17'b10101011101000000;
uRam[734 ] <= 17'b10101011111000000;
uRam[735 ] <= 17'b01100001100100001;
uRam[736 ] <= 17'b00000000000000000;
uRam[737 ] <= 17'b00000000000000000;
uRam[738 ] <= 17'b00000000000000000;
uRam[739 ] <= 17'b00000000000000000;
uRam[740 ] <= 17'b00000000000000000;
uRam[741 ] <= 17'b00000000000000000;
uRam[742 ] <= 17'b00000000000000000;
uRam[743 ] <= 17'b00000000000000000;
uRam[744 ] <= 17'b00000000000000000;
uRam[745 ] <= 17'b00000000000000000;
uRam[746 ] <= 17'b00000000000000000;
uRam[747 ] <= 17'b00000000000000000;
uRam[748 ] <= 17'b00000000000000000;
uRam[749 ] <= 17'b00000000000000000;
uRam[750 ] <= 17'b00000000000000000;
uRam[751 ] <= 17'b00000000000000000;
uRam[752 ] <= 17'b00110010100111010;
uRam[753 ] <= 17'b10001010010100001;
uRam[754 ] <= 17'b10110100100000000;
uRam[755 ] <= 17'b10110100111000001;
uRam[756 ] <= 17'b01110010110111010;
uRam[757 ] <= 17'b10001010010100001;
uRam[758 ] <= 17'b10101011010100000;
uRam[759 ] <= 17'b10110100110100001;
uRam[760 ] <= 17'b10111100100100001;
uRam[761 ] <= 17'b01101111110000000;
uRam[762 ] <= 17'b01000110010000001;
uRam[763 ] <= 17'b10101111111100000;
uRam[764 ] <= 17'b10101011110000001;
uRam[765 ] <= 17'b01100011110000000;
uRam[766 ] <= 17'b01110100100100001;
uRam[767 ] <= 17'b10110000000000000;
uRam[768 ] <= 17'b10011001110000000;
uRam[769 ] <= 17'b00110110000000000;
uRam[770 ] <= 17'b00101111001000000;
uRam[771 ] <= 17'b10111110000100000;
uRam[772 ] <= 17'b00110100111000000;
uRam[773 ] <= 17'b10001100100100000;
uRam[774 ] <= 17'b00000000000000100;
uRam[775 ] <= 17'b00110010000000000;
uRam[776 ] <= 17'b00000100010100110;
uRam[777 ] <= 17'b00111110000100000;
uRam[778 ] <= 17'b00111110000100000;
uRam[779 ] <= 17'b10100111011000000;
uRam[780 ] <= 17'b01110100110000001;
uRam[781 ] <= 17'b01110100100100000;
uRam[782 ] <= 17'b10010101000000000;
uRam[783 ] <= 17'b10110110100000000;
uRam[784 ] <= 17'b00000000000000000;
uRam[785 ] <= 17'b00000000000000000;
uRam[786 ] <= 17'b00000000000000000;
uRam[787 ] <= 17'b00000000000000000;
uRam[788 ] <= 17'b00000000000000000;
uRam[789 ] <= 17'b00000000000000000;
uRam[790 ] <= 17'b00000000000000000;
uRam[791 ] <= 17'b00000000000000000;
uRam[792 ] <= 17'b00000000000000000;
uRam[793 ] <= 17'b00000000000000000;
uRam[794 ] <= 17'b00000000000000000;
uRam[795 ] <= 17'b00000000000000000;
uRam[796 ] <= 17'b00000000000000000;
uRam[797 ] <= 17'b00000000000000000;
uRam[798 ] <= 17'b00000000000000000;
uRam[799 ] <= 17'b00000000000000000;
uRam[800 ] <= 17'b00110110000000000;
uRam[801 ] <= 17'b00010110001100000;
uRam[802 ] <= 17'b00000110010111010;
uRam[803 ] <= 17'b00000110010111010;
uRam[804 ] <= 17'b00110100111000000;
uRam[805 ] <= 17'b10111010010000000;
uRam[806 ] <= 17'b00001110110000000;
uRam[807 ] <= 17'b00000000000000100;
uRam[808 ] <= 17'b10110000110100001;
uRam[809 ] <= 17'b01111010100000000;
uRam[810 ] <= 17'b01010110001100001;
uRam[811 ] <= 17'b10111010110000000;
uRam[812 ] <= 17'b10110000110100000;
uRam[813 ] <= 17'b00100001010001010;
uRam[814 ] <= 17'b01010110001100001;
uRam[815 ] <= 17'b01110000100100000;
uRam[816 ] <= 17'b00000000000000000;
uRam[817 ] <= 17'b00000000000000000;
uRam[818 ] <= 17'b00000000000000000;
uRam[819 ] <= 17'b00000000000000000;
uRam[820 ] <= 17'b00000000000000000;
uRam[821 ] <= 17'b00000000000000000;
uRam[822 ] <= 17'b00000000000000000;
uRam[823 ] <= 17'b00000000000000000;
uRam[824 ] <= 17'b00000000000000000;
uRam[825 ] <= 17'b00000000000000000;
uRam[826 ] <= 17'b00000000000000000;
uRam[827 ] <= 17'b00000000000000000;
uRam[828 ] <= 17'b00000000000000000;
uRam[829 ] <= 17'b00000000000000000;
uRam[830 ] <= 17'b00000000000000000;
uRam[831 ] <= 17'b00000000000000000;
uRam[832 ] <= 17'b00000100111000000;
uRam[833 ] <= 17'b10111000000100001;
uRam[834 ] <= 17'b00000000000000100;
uRam[835 ] <= 17'b00110000010100000;
uRam[836 ] <= 17'b01111110000100000;
uRam[837 ] <= 17'b10111000010100001;
uRam[838 ] <= 17'b00000000000000100;
uRam[839 ] <= 17'b00111000001100000;
uRam[840 ] <= 17'b01111110000100000;
uRam[841 ] <= 17'b10000000000000100;
uRam[842 ] <= 17'b01111100100100000;
uRam[843 ] <= 17'b01000000000000100;
uRam[844 ] <= 17'b00000000000000100;
uRam[845 ] <= 17'b01110100111000000;
uRam[846 ] <= 17'b01111100110100000;
uRam[847 ] <= 17'b01110010100100000;
uRam[848 ] <= 17'b00000000000000000;
uRam[849 ] <= 17'b00000000000000000;
uRam[850 ] <= 17'b00000000000000000;
uRam[851 ] <= 17'b00000000000000000;
uRam[852 ] <= 17'b00000000000000000;
uRam[853 ] <= 17'b00000000000000000;
uRam[854 ] <= 17'b00000000000000000;
uRam[855 ] <= 17'b00000000000000000;
uRam[856 ] <= 17'b00000000000000000;
uRam[857 ] <= 17'b00000000000000000;
uRam[858 ] <= 17'b00000000000000000;
uRam[859 ] <= 17'b00000000000000000;
uRam[860 ] <= 17'b00000000000000000;
uRam[861 ] <= 17'b00000000000000000;
uRam[862 ] <= 17'b00000000000000000;
uRam[863 ] <= 17'b00000000000000000;
uRam[864 ] <= 17'b01001110111100000;
uRam[865 ] <= 17'b00000000000000100;
uRam[866 ] <= 17'b00000000000000100;
uRam[867 ] <= 17'b10110000110100001;
uRam[868 ] <= 17'b00000000000000000;
uRam[869 ] <= 17'b00000000000000000;
uRam[870 ] <= 17'b00000000000000000;
uRam[871 ] <= 17'b01011001100000000;
uRam[872 ] <= 17'b01111010100100001;
uRam[873 ] <= 17'b00000000001001010;
uRam[874 ] <= 17'b10000000000000100;
uRam[875 ] <= 17'b01110010110100000;
uRam[876 ] <= 17'b01110110110100000;
uRam[877 ] <= 17'b01111010110100001;
uRam[878 ] <= 17'b01111110000100000;
uRam[879 ] <= 17'b00000000000000100;
uRam[880 ] <= 17'b00000000000000000;
uRam[881 ] <= 17'b00000000000000000;
uRam[882 ] <= 17'b00000000000000000;
uRam[883 ] <= 17'b00000000000000000;
uRam[884 ] <= 17'b00000000000000000;
uRam[885 ] <= 17'b00000000000000000;
uRam[886 ] <= 17'b00000000000000000;
uRam[887 ] <= 17'b00000000000000000;
uRam[888 ] <= 17'b00000000000000000;
uRam[889 ] <= 17'b00000000000000000;
uRam[890 ] <= 17'b00000000000000000;
uRam[891 ] <= 17'b00000000000000000;
uRam[892 ] <= 17'b00000000000000000;
uRam[893 ] <= 17'b00000000000000000;
uRam[894 ] <= 17'b00000000000000000;
uRam[895 ] <= 17'b00000000000000000;
uRam[896 ] <= 17'b10001100110100111;
uRam[897 ] <= 17'b10111100001000001;
uRam[898 ] <= 17'b10111100001000001;
uRam[899 ] <= 17'b00101101000000110;
uRam[900 ] <= 17'b10001100101100111;
uRam[901 ] <= 17'b10111100011000001;
uRam[902 ] <= 17'b10111100011000001;
uRam[903 ] <= 17'b00101101010000110;
uRam[904 ] <= 17'b10110100101000000;
uRam[905 ] <= 17'b01111110000100000;
uRam[906 ] <= 17'b10110100101000000;
uRam[907 ] <= 17'b10111100100100001;
uRam[908 ] <= 17'b10111110110000000;
uRam[909 ] <= 17'b01000000000000100;
uRam[910 ] <= 17'b10111110110000000;
uRam[911 ] <= 17'b10111000100100001;
uRam[912 ] <= 17'b00000000000000000;
uRam[913 ] <= 17'b00000000000000000;
uRam[914 ] <= 17'b00000000000000000;
uRam[915 ] <= 17'b00000000000000000;
uRam[916 ] <= 17'b00000000000000000;
uRam[917 ] <= 17'b00000000000000000;
uRam[918 ] <= 17'b00000000000000000;
uRam[919 ] <= 17'b00000000000000000;
uRam[920 ] <= 17'b00000000000000000;
uRam[921 ] <= 17'b00000000000000000;
uRam[922 ] <= 17'b00000000000000000;
uRam[923 ] <= 17'b00000000000000000;
uRam[924 ] <= 17'b00000000000000000;
uRam[925 ] <= 17'b00000000000000000;
uRam[926 ] <= 17'b00000000000000000;
uRam[927 ] <= 17'b00000000000000000;
uRam[928 ] <= 17'b10111110000000000;
uRam[929 ] <= 17'b10110010010000001;
uRam[930 ] <= 17'b00111110010000001;
uRam[931 ] <= 17'b00111000001100000;
uRam[932 ] <= 17'b10101001110000000;
uRam[933 ] <= 17'b10110000000100001;
uRam[934 ] <= 17'b00101111100100000;
uRam[935 ] <= 17'b00111000101110000;
uRam[936 ] <= 17'b00110010100111010;
uRam[937 ] <= 17'b01111010101000000;
uRam[938 ] <= 17'b01000110010000001;
uRam[939 ] <= 17'b01000110010000000;
uRam[940 ] <= 17'b01110010110111010;
uRam[941 ] <= 17'b01111010111000000;
uRam[942 ] <= 17'b01110100100100001;
uRam[943 ] <= 17'b01110100100100001;
uRam[944 ] <= 17'b00000000000000000;
uRam[945 ] <= 17'b00000000000000000;
uRam[946 ] <= 17'b00000000000000000;
uRam[947 ] <= 17'b00000000000000000;
uRam[948 ] <= 17'b00000000000000000;
uRam[949 ] <= 17'b00000000000000000;
uRam[950 ] <= 17'b00000000000000000;
uRam[951 ] <= 17'b00000000000000000;
uRam[952 ] <= 17'b00000000000000000;
uRam[953 ] <= 17'b00000000000000000;
uRam[954 ] <= 17'b00000000000000000;
uRam[955 ] <= 17'b00000000000000000;
uRam[956 ] <= 17'b00000000000000000;
uRam[957 ] <= 17'b00000000000000000;
uRam[958 ] <= 17'b00000000000000000;
uRam[959 ] <= 17'b00000000000000000;
uRam[960 ] <= 17'b00101001110100000;
uRam[961 ] <= 17'b10001100100100000;
uRam[962 ] <= 17'b01110010000100000;
uRam[963 ] <= 17'b10110000110100001;
uRam[964 ] <= 17'b00000010000011110;
uRam[965 ] <= 17'b01111000000000000;
uRam[966 ] <= 17'b01000000101000000;
uRam[967 ] <= 17'b10110000010000001;
uRam[968 ] <= 17'b00101101110100000;
uRam[969 ] <= 17'b10111010000000000;
uRam[970 ] <= 17'b01001010001000000;
uRam[971 ] <= 17'b10110110000100001;
uRam[972 ] <= 17'b00000000000000000;
uRam[973 ] <= 17'b00000000000000000;
uRam[974 ] <= 17'b00000000000000000;
uRam[975 ] <= 17'b00000000000000000;
uRam[976 ] <= 17'b00000000000000000;
uRam[977 ] <= 17'b00000000000000000;
uRam[978 ] <= 17'b00000000000000000;
uRam[979 ] <= 17'b00000000000000000;
uRam[980 ] <= 17'b00000000000000000;
uRam[981 ] <= 17'b00000000000000000;
uRam[982 ] <= 17'b00000000000000000;
uRam[983 ] <= 17'b00000000000000000;
uRam[984 ] <= 17'b00000000000000000;
uRam[985 ] <= 17'b00000000000000000;
uRam[986 ] <= 17'b00000000000000000;
uRam[987 ] <= 17'b00000000000000000;
uRam[988 ] <= 17'b00000000000000000;
uRam[989 ] <= 17'b00000000000000000;
uRam[990 ] <= 17'b00000000000000000;
uRam[991 ] <= 17'b00000000000000000;
uRam[992 ] <= 17'b10100111101000000;
uRam[993 ] <= 17'b00000000000000000;
uRam[994 ] <= 17'b10010010000000010;
uRam[995 ] <= 17'b10100111000000001;
uRam[996 ] <= 17'b10100111111000000;
uRam[997 ] <= 17'b00000000000000000;
uRam[998 ] <= 17'b10010010010000010;
uRam[999 ] <= 17'b10001110011100001;
uRam[1000] <= 17'b00100011001100000;
uRam[1001] <= 17'b00100001001001010;
uRam[1002] <= 17'b10010011000000010;
uRam[1003] <= 17'b10001010110100001;
uRam[1004] <= 17'b01100011011100000;
uRam[1005] <= 17'b00100001011001010;
uRam[1006] <= 17'b10010011010000010;
uRam[1007] <= 17'b10001010100100001;
uRam[1008] <= 17'b00000000000000000;
uRam[1009] <= 17'b00000000000000000;
uRam[1010] <= 17'b00000000000000000;
uRam[1011] <= 17'b00000000000000000;
uRam[1012] <= 17'b00000000000000000;
uRam[1013] <= 17'b00000000000000000;
uRam[1014] <= 17'b00000000000000000;
uRam[1015] <= 17'b00000000000000000;
uRam[1016] <= 17'b00000000000000000;
uRam[1017] <= 17'b00000000000000000;
uRam[1018] <= 17'b00000000000000000;
uRam[1019] <= 17'b00000000000000000;
uRam[1020] <= 17'b00000000000000000;
uRam[1021] <= 17'b00000000000000000;
uRam[1022] <= 17'b00000000000000000;
uRam[1023] <= 17'b00000000000000000;

	end
	
	always @( posedge clk) microOutput <= uRam[ microAddr];
endmodule


module nanoRom( input clk, input [NADDR_WIDTH-1:0] nanoAddr, output reg [NANO_WIDTH-1:0] nanoOutput);
	reg [NANO_WIDTH-1:0] nRam[ NANO_DEPTH];		
	initial begin
nRam[0  ] <= 68'b00000000000000000000000000000000000000000000000010000000000000000000;
nRam[1  ] <= 68'b00000000000000000000000000000000000000000000000010000000000000000000;
nRam[2  ] <= 68'b00000000000000000000000000000000000000000000000010000000000000000000;
nRam[3  ] <= 68'b00000000000000000000000000001000000110011100000000000000101001000001;
nRam[4  ] <= 68'b00100001000000011000010001001000000110100000000001000000011001001001;
nRam[5  ] <= 68'b00000001100000000010100000001000000110000000001001000000001001001001;
nRam[6  ] <= 68'b00100000000000011000010001000000000101000000000010000000100001010000;
nRam[7  ] <= 68'b11000001000000000000000000001000000100010000000001000000000001010001;
nRam[8  ] <= 68'b00100001000000011000010000000000000000000000000101000000000000010000;
nRam[9  ] <= 68'b01000001011000000000100000000110010001000000001100000000110100011000;
nRam[10 ] <= 68'b01000001011000000000100000000110010001000000001100000001100100011000;
nRam[11 ] <= 68'b00100001000000011000010000000000000100000000000001000000000001010000;
nRam[12 ] <= 68'b10100100001000011000001000010000101001110000000001000100110010100001;
nRam[13 ] <= 68'b01000000000000000000000010000000010100000000001000110001000000000000;
nRam[14 ] <= 68'b00100001000000011000000000110010100100011111010001100000000001000000;
nRam[15 ] <= 68'b00100010000000011000000000000000100010000100000000010100000100000011;
nRam[16 ] <= 68'b00000001011000000000000001000110000000000000000010000000000100000000;
nRam[17 ] <= 68'b00000000000000000000000000001000000100000000000001000000000001010001;
nRam[18 ] <= 68'b00000001100000000010100000001000000110000000001001010000001001001001;
nRam[19 ] <= 68'b00101000000000001000010000000000000000000000000010000000000000000000;
nRam[20 ] <= 68'b01100010000000011000010010000000010100000000001000110001000000000000;
nRam[21 ] <= 68'b00000000000000000000000010010010100000000000000100110010000000000000;
nRam[22 ] <= 68'b00100000000000011000010001001000000110000000001001010000001001001001;
nRam[23 ] <= 68'b00000000000000000000001000000000100100000000000000110010000001011000;
nRam[24 ] <= 68'b00010010000000000100100000001000000100000000000010000000000001010001;
nRam[25 ] <= 68'b00100010000000011100000000000000000001100000000010001000100000000000;
nRam[26 ] <= 68'b00010010000000000100000000000000010001100000000010000000000000000000;
nRam[27 ] <= 68'b00000000000000000000000000011001100110100000010001000000011011010001;
nRam[28 ] <= 68'b10100010110000000000000000000000100000010000010010000100000100000000;
nRam[29 ] <= 68'b10000000000000000000000000001000000100010000000001000000000001000001;
nRam[30 ] <= 68'b00100000000000011001000000011010000110000000001001000000001001001001;
nRam[31 ] <= 68'b00010011000000000000101000010000001001000000010101000000100000110000;
nRam[32 ] <= 68'b00000001000000000001010000000000000000000000000101100000000000010000;
nRam[33 ] <= 68'b00100010000000011000001000001000100110000000000001000000000001010001;
nRam[34 ] <= 68'b00000001000000000010100001010000001001000000010110000000100000110000;
nRam[35 ] <= 68'b01000001000000000000000000000000000001101010001100000000110000000000;
nRam[36 ] <= 68'b00110100000000000100000100000000000000000000000010000000000000000000;
nRam[37 ] <= 68'b00000000000100100000100000000000010000000000000000000001000000011000;
nRam[38 ] <= 68'b01110101000000000100100000100010000001100000000000000000110100001010;
nRam[39 ] <= 68'b00100010000000011010000100000000100010000100000000010100000100000011;
nRam[40 ] <= 68'b11000001000000000000000000001000000100010000000001000000000001010001;
nRam[41 ] <= 68'b01010011000000000100100000100010000001100000000000000000110100001010;
nRam[42 ] <= 68'b11000001000000000000000000001001100110110000000001000000011011000001;
nRam[43 ] <= 68'b01001001110000000000001000001000001000000000000101000000000000100001;
nRam[44 ] <= 68'b00000000000000000000100000100010010000000000000000110001000100000010;
nRam[45 ] <= 68'b00010000110000000001010000000000000000011100000010000000000000011000;
nRam[46 ] <= 68'b01010001110000000001000000011010100100000000000001000000000001000001;
nRam[47 ] <= 68'b00000000000000000000000001000000000100000000001100010000000001010000;
nRam[48 ] <= 68'b00001000000000011001001000001000000110100000000001000100000011010001;
nRam[49 ] <= 68'b01010001110000000001010000001000001000000000000101000000000000110001;
nRam[50 ] <= 68'b10100010110100100100000001000000000001110000000010000000110000010000;
nRam[51 ] <= 68'b00000000000100000000000000000010100001001010000101100000100000010000;
nRam[52 ] <= 68'b00010000110000000001000000000000100000000000010010000100000100000000;
nRam[53 ] <= 68'b10000000000000000000000000001000000100010000000001000000000001000001;
nRam[54 ] <= 68'b00000001000000000000000001000000001001000000000101000000100000100000;
nRam[55 ] <= 68'b00010010000000000000100000001010101000000000000101000000000000110001;
nRam[56 ] <= 68'b10100000000100111000000000100001100010111010000101100000011010010010;
nRam[57 ] <= 68'b00100000000000011000000000110010100110000000010000100000001101000010;
nRam[58 ] <= 68'b00010010000000001100000000000000000000000000000010000000000000000000;
nRam[59 ] <= 68'b11000001000000000000001000011101100100010000000001000000000001000001;
nRam[60 ] <= 68'b00010100000000000100000100000000000000000000000010000000000000000000;
nRam[61 ] <= 68'b10100010110000000100001000000000100000010000010010000100000010000000;
nRam[62 ] <= 68'b00100000000100111000000000000000100000010010000101000100000100010010;
nRam[63 ] <= 68'b00100010000000011000000000000000100010000100000000010100000100000011;
nRam[64 ] <= 68'b00100010100000011001010000010000100100000000001110000100001000000000;
nRam[65 ] <= 68'b00000000000100000000000000000010100000001010000101000000000000010000;
nRam[66 ] <= 68'b00100010100000011001000000010010100100000000001110000100001000000000;
nRam[67 ] <= 68'b00000001000000000000010000000000100000000000010101000100000010010000;
nRam[68 ] <= 68'b00000000000100100000000000100010000000000100000000110001000100011010;
nRam[69 ] <= 68'b00100000000000011000000000010000100110000000011000100000001001000000;
nRam[70 ] <= 68'b00000000000100100000100000100010010000000000000000110001000100011010;
nRam[71 ] <= 68'b00000000011000000000000000000110000000000000001110000000110100111000;
nRam[72 ] <= 68'b00011000000000011001001000001000000100000000000001000000000001010001;
nRam[73 ] <= 68'b00100010000000011100000000000000000001100000000010001000100000000000;
nRam[74 ] <= 68'b00110000100000001000000100000000100000000000000010000100000100000000;
nRam[75 ] <= 68'b00000000000100000000000000000010100001000000000101100000100000010000;
nRam[76 ] <= 68'b10100010110000000100001000010001100000010000000010000000000000000000;
nRam[77 ] <= 68'b01000001000000000000000000000000000000000000000101000000000000010000;
nRam[78 ] <= 68'b10000000000000000000000000001000000100010000000001000000000001000001;
nRam[79 ] <= 68'b00000000000000000000000000001000001000000000000101000000000000110001;
nRam[80 ] <= 68'b00001000110000000000001000000000000000000000000010000000000000000000;
nRam[81 ] <= 68'b00010010000000001100000000000000000000000000000010000000000000000000;
nRam[82 ] <= 68'b00010000000000001010000100000000110001000000000010000100011000000000;
nRam[83 ] <= 68'b01010001000000011000001000000000000001100000000000000000110000000000;
nRam[84 ] <= 68'b00001100000000011000001000100001000010100000000101110000000000000011;
nRam[85 ] <= 68'b01000000000000000000000010000000010100000000001000110000000001000000;
nRam[86 ] <= 68'b11000001000000000000000000001000001000010000000101000000000000100001;
nRam[87 ] <= 68'b00000000000000000000000000001000000100011100000001100000000001000001;
nRam[88 ] <= 68'b00000000000000000000000000000000000000000000000101100000000000000000;
nRam[89 ] <= 68'b00000000000100000000000000000000100000000000000101000100000100010000;
nRam[90 ] <= 68'b11101011000000000000000000000000000000010000000010000000000000000000;
nRam[91 ] <= 68'b01100001000000011001000000011010100100000000000001000000000001000001;
nRam[92 ] <= 68'b01100010000000011000010010000000010100000000001000110000000001000000;
nRam[93 ] <= 68'b00000000000000000000000010010010100000000000010100110000000100000000;
nRam[94 ] <= 68'b01000001000000000000010000011001101000000000000101000100001000110001;
nRam[95 ] <= 68'b00100000000100111100000000000000000010000010000100100010001000010000;
nRam[96 ] <= 68'b00010010000000000000000000000010110100000000001110000000000000011000;
nRam[97 ] <= 68'b00000000000000000000001000010000100100000000011100110010000001011000;
nRam[98 ] <= 68'b00000000000100000000000000010000111000000000010101000100011000110000;
nRam[99 ] <= 68'b00000000011000000010100000000110000100000000001101110000000101000000;
nRam[100] <= 68'b00000000000000000000000000000000000000000000000010000000000000000000;
nRam[101] <= 68'b00000001000000000000000000000000010101001010001101000000100001010000;
nRam[102] <= 68'b00000001000000000000010000000000100000000000000101000100001000010000;
nRam[103] <= 68'b01110101000000010000001000000000000001100000000000000000110000000000;
nRam[104] <= 68'b01000001000000000000000010000000010100001010001000110001000000000000;
nRam[105] <= 68'b00100010000000011000000000011010101010000000010101000000001100110001;
nRam[106] <= 68'b00100001000000011000010001010000000100000000010000010000000001010000;
nRam[107] <= 68'b01000001000000000000010000000000100000000110000101000000000000010000;
nRam[108] <= 68'b01000001000000000000000010000000010100001010001000110001000000000000;
nRam[109] <= 68'b00100000000000011000010001010001000000000000011010000000000010001000;
nRam[110] <= 68'b00000001000000000000000001010000000100000000010001110000000001000000;
nRam[111] <= 68'b00010010000000001000000000011010101000000000000101000000000000110001;
nRam[112] <= 68'b00000000000000000000000000001000001000000000000101000000000000110001;
nRam[113] <= 68'b00010010000000000001100000000010000000000000000101100000000000000000;
nRam[114] <= 68'b00010010000000000001000000000010000100000000000101100000000000000000;
nRam[115] <= 68'b00100010000000011100000000001000001000000000000101000000000000100001;
nRam[116] <= 68'b00000001000000000001010000000000001010100000000110000000011000101000;
nRam[117] <= 68'b00000001100000000000100000000000000000000000000101000000000000010000;
nRam[118] <= 68'b00010010000000000000101000001001000100000000001001000000000011010001;
nRam[119] <= 68'b11110101001000000100000000000000000000010000000010000000000000000000;
nRam[120] <= 68'b00000000000000000000010000001001101000000000000101000010000010110001;
nRam[121] <= 68'b00000000000000000000010000000000100000000110000101100000000000000000;
nRam[122] <= 68'b00100010100000001001100000000010000010000100001000000000001000001000;
nRam[123] <= 68'b00100010100000001001000000000010000110000100001000000000001000001000;
nRam[124] <= 68'b00010010000000001000010000000000000000000000001110000000000000011000;
nRam[125] <= 68'b00110100000100101100000000000000000001100000000001100000110000010000;
nRam[126] <= 68'b01110101000000001000000100000000111000000000010010000100000100000000;
nRam[127] <= 68'b01000000000000000000010000010000100110000000011100100000000001011000;
nRam[128] <= 68'b11010011000000000000101000001001000100010000001001000000000011010001;
nRam[129] <= 68'b11110101001000000000000000000000100000010000000010000100000100000000;
nRam[130] <= 68'b01110101000000000100000000000000010000000000010010001000000001000000;
nRam[131] <= 68'b01110101000000000000000000000000110000000000010010001100000101000000;
nRam[132] <= 68'b01110101000000000000000000000000110000000000010010001100011001000000;
nRam[133] <= 68'b01110000000000011100000000000000000001100000001101000000110000000000;
nRam[134] <= 68'b00010000000000001000000000000010100000000000000010000000000000000000;
nRam[135] <= 68'b00010010000000000100000100000000010001000000000010000000000000000000;
nRam[136] <= 68'b01000000000000000000010000010000100110000000011100100010001001011000;
nRam[137] <= 68'b00100000000000011000010000000000000100000000000000100000000001000000;
nRam[138] <= 68'b00000001000000000000000000000000001000000000000101000000000000110000;
nRam[139] <= 68'b00100001000000011100000001011001000110000000011000000000001011001001;
nRam[140] <= 68'b01100001000000011000000000010010100110000000011100100000001101011000;
nRam[141] <= 68'b01100001000000011000010000010010000010000000010101000000001100010000;
nRam[142] <= 68'b00000000000000000000000100000000010010100000001100110001011000011000;
nRam[143] <= 68'b01100001000000011000000000010000100110000000011000100000001001000000;
nRam[144] <= 68'b00000000000000000000000000001000000100011100000001100000000001000001;
nRam[145] <= 68'b00010010000000000000000000010010110110000000001110000010001000011000;
nRam[146] <= 68'b01000001000000000000100000010010010000000000010000110001000100011000;
nRam[147] <= 68'b00010010000000000000010000010000110110000000001110000010001000011000;
nRam[148] <= 68'b01000001000000000000000010000000010100001010001000110000000001000000;
nRam[149] <= 68'b01000001000000000000010000001000101000000110000101000000000000110001;
nRam[150] <= 68'b00000001000000000000010000000000100000000000000101000100001000010000;
nRam[151] <= 68'b00101000000000001000010000000000000000000000000010000000000000000000;
nRam[152] <= 68'b00100010000000011000000000000000100000000000000010000100011000000000;
nRam[153] <= 68'b00100010001000011010000000000000100000000000000010000100000100000000;
nRam[154] <= 68'b11010011001000000100000000010000011000010000000010000000000000000000;
nRam[155] <= 68'b00010010000000000100000000000000010000000000010010001000000001000000;
nRam[156] <= 68'b00001000000000011000001000000000000000000000000101110000000000000011;
nRam[157] <= 68'b00100010110000000000010000001000001000000000000101000000000000110001;
nRam[158] <= 68'b00100010000000011000000000000000100010100000000010000000000000000000;
nRam[159] <= 68'b00100000000000011000000000110001100100011111011001100000000011000010;
nRam[160] <= 68'b00100000000000011000000000001000100110000000001001010000001001000001;
nRam[161] <= 68'b01000001000000000000000000010000000100000000011100100000000001011000;
nRam[162] <= 68'b00000000100000000010100000000000000001000000000101000000100000010000;
nRam[163] <= 68'b00000001000000000000000000011001000100000000011001000000000011000001;
nRam[164] <= 68'b00000000011000000010100001000110000101000000000000010000100101010000;
nRam[165] <= 68'b00100001000000011100000001011001000100000000011001000000000011000001;
nRam[166] <= 68'b01000000000000000000000000000000000101001010001101100000100001000000;
nRam[167] <= 68'b00000000000100000000000000000000100001001010000101100100100100010000;
nRam[168] <= 68'b00000000011000000000000000000010110110000000001100000000001101011000;
nRam[169] <= 68'b01000001000000000000000000000001111001100000001010000000110010100000;
nRam[170] <= 68'b00110010000000011000000000010010100010000000001110000010001000011000;
nRam[171] <= 68'b11000001000000000000000000011001100110110000010001000000011011000001;
nRam[172] <= 68'b00100000000000011010000000100001110000001100001010000000000010000010;
nRam[173] <= 68'b00000000000000000000000000010000000100010101010001100000000001000000;
nRam[174] <= 68'b01000000000000000000000000000000000010100000000010000000011000001000;
nRam[175] <= 68'b00000001000000000000000000000000000001101010001101000000110000010000;
nRam[176] <= 68'b10000000000000000000001000001101100100010000000001000000000001000001;
nRam[177] <= 68'b01110101000000000000000000000000110000000000000010001100000101000000;
nRam[178] <= 68'b11000001000000000000000000001000000100010000000001000000000001000001;
nRam[179] <= 68'b00100010000000011000000000001001101000000010000101000010000010110001;
nRam[180] <= 68'b00100010000100011000000000010010100000000000000101000000000000010000;
nRam[181] <= 68'b11100101000000011100000000001001000100010000001001000000000011010001;
nRam[182] <= 68'b00100100000100111000000000000000100000000000010101100100000100010000;
nRam[183] <= 68'b00100010000100011000000000011010100100000000000000000000000001011001;
nRam[184] <= 68'b00100000000000001000001000000000100000000000000010000100000010000000;
nRam[185] <= 68'b00100010000000011100001000001000100100000000000001000100001001010001;
nRam[186] <= 68'b00010010000000000100000100000000010001000000000010000000000000000000;
nRam[187] <= 68'b10000000000000000000001000011101000100010000000001000000000001000001;
nRam[188] <= 68'b00011000000000011000001000000000100010000000000010000000000000000000;
nRam[189] <= 68'b01000000000000000000000000000000000100000000000001000000000001010000;
nRam[190] <= 68'b01000000000000000000010000010000100110000000011100100000011001001000;
nRam[191] <= 68'b00000000001000000010001000010001010000000000000010001000000000100000;
nRam[192] <= 68'b11100101000000011100000000001000001000010000000101000000000000110001;
nRam[193] <= 68'b01000001000000000000001000010001100000000000000010000000000000000000;
nRam[194] <= 68'b00110100000000000000000000000000110000000000000010001100000101000000;
nRam[195] <= 68'b10000000000000000000001000001000100100010000010001000100000011000001;
nRam[196] <= 68'b01110101000000000100001000000001110000000000010010001000000001000000;
nRam[197] <= 68'b10000000000000000000001000001000100100010000000001000100000011000001;
nRam[198] <= 68'b00110100000000000000000000000000110000000000010010001100000101000000;
nRam[199] <= 68'b00110100000000000000000000000000110000000000010010001100011001000000;
nRam[200] <= 68'b01000000000000000000000000010000000110100000011100100000011001001000;
nRam[201] <= 68'b00000000000100000000000000010000111000000000010101000100000100110010;
nRam[202] <= 68'b00000000000100000000000000100010100001100000000001000000110000011000;
nRam[203] <= 68'b01000000000000000000000000010010000110000000010000100000001101001000;
nRam[204] <= 68'b00000000000000000000000000001000000110000000001001000000001001001001;
nRam[205] <= 68'b01000000000000000000010000000001100000000000000101000010000010010000;
nRam[206] <= 68'b01000000000000000000000000001000000110000000001001010000001001000001;
nRam[207] <= 68'b00000001000000000000000000000000000001101010001101000000110000000000;
nRam[208] <= 68'b11100101000000011000000000010000111001110000010010000100110100100000;
nRam[209] <= 68'b00000000000000000000000000011010101010000000000101000010001000110001;
nRam[210] <= 68'b11000001000000000000001000001101100100010000000001000000000001000001;
nRam[211] <= 68'b00000000000000000000000100000000010000000000000001100001000000000000;
nRam[212] <= 68'b00000000000000000000000000001001100100000000001001000000000011010001;
nRam[213] <= 68'b11000001000000000000010000010001100000010000010010000000011010000000;
nRam[214] <= 68'b00000000000000000000000000000000000000010110000010000000000000000000;
nRam[215] <= 68'b00000000000000000000000000000000000000001100000000000001000000000000;
nRam[216] <= 68'b00100010000000011000000000000000100010100000000010000000000000000000;
nRam[217] <= 68'b00001000000000011000001000000000000000000000000101110000000000000011;
nRam[218] <= 68'b10000000000000000000000000000000000000010000000010000000000000000000;
nRam[219] <= 68'b00000000000000000000010000000000100010000000000010000010001000000000;
nRam[220] <= 68'b00101000000000001000001000000000000000000000000010000000000000000000;
nRam[221] <= 68'b01010011000000000000100000000010100001100000001100000000110000011000;
nRam[222] <= 68'b00000001000010000000000001000000000000000000000101000000000000010000;
nRam[223] <= 68'b00100010000000011000010000001101101000000000000101000000000000110001;
nRam[224] <= 68'b00000000000000000000100000010010010000000000010000110001000100000000;
nRam[225] <= 68'b01000000000000000000000000010000000100000000011100100000000001000000;
nRam[226] <= 68'b00000000000000000000000100010010010000000000010000110001000100000000;
nRam[227] <= 68'b01000000000000000000100000000000010000000000000001000000110000010000;
nRam[228] <= 68'b01010011000000001000010000000000000001100000001100000000110000011000;
nRam[229] <= 68'b01000001000000000000010000001001101000000000000101000000000000110001;
nRam[230] <= 68'b00100100000100011001000000000000100000000000010101000100000100010000;
nRam[231] <= 68'b01100010000000011000100000010010110010000000001100000000110000011000;
nRam[232] <= 68'b00011000000000011000001000000000000000000000000101110000000000000011;
nRam[233] <= 68'b00000000000000000000000000001000000100000000000001000000000001010001;
nRam[234] <= 68'b00010010000000000100000100000000010001000000000010000000000000000000;
nRam[235] <= 68'b00001010000000011000001000000000000000000000000101110000000000000011;
nRam[236] <= 68'b00010010000000000000000000000001110100000010001110000010000010011000;
nRam[237] <= 68'b01100010000000011000100000010010110010000000001100000001000000011000;
nRam[238] <= 68'b01000000000000000000100000000010010000000000001100110001000100011000;
nRam[239] <= 68'b00100010000100011000000001011010100100000000000001000000000001011001;
nRam[240] <= 68'b00000001000000000000010000000001100001001010000101000000100000010000;
nRam[241] <= 68'b00000000000000000000010000000000100101000110001110000000100001011000;
nRam[242] <= 68'b00000000000000000000100000010010010000000000010000110001000100011000;
nRam[243] <= 68'b01010011000000000000100000000001100001100010001100000010110010011000;
nRam[244] <= 68'b01100011000000011000000000010010100100000000011101110000000001011000;
nRam[245] <= 68'b00000000000100000001000000010000100100000000011101000100000101010000;
nRam[246] <= 68'b00100010000100011000000001010010100100000000011100010000000001010000;
nRam[247] <= 68'b00000001000000000000010000000000100000000001000101000100000010010000;
nRam[248] <= 68'b00000001000000000000010000000001100000001111000101000000000000010000;
nRam[249] <= 68'b00000000000000000000000000010010100000000110010101100000000100000000;
nRam[250] <= 68'b00000111000000000000010000010000111000001000010110000100001000100000;
nRam[251] <= 68'b01000000000000000000100000000001110000000000001001000000110010010000;
nRam[252] <= 68'b01001011000000011000001000000000000001100000000000000000110000000000;
nRam[253] <= 68'b00000000000000000000010000000000100010000000000101000000000000010000;
nRam[254] <= 68'b10100100000000011100000000001000000100010000000001000000000001000001;
nRam[255] <= 68'b00010000000000000000000000010000100100000010000010000000000000000000;
nRam[256] <= 68'b00000000000000000000000000001000000100000010000000110010000001000001;
nRam[257] <= 68'b01000000000000000000000000001001100100000000001001010000000011000001;
nRam[258] <= 68'b00000000000000000000000000001001100100000000001001010000000011000001;
nRam[259] <= 68'b00100000000000011000000000010010100010000000010101000000001100010000;
nRam[260] <= 68'b00000000000100000000000000000000101000000000000101000100011000110000;
nRam[261] <= 68'b00000000000100100000100000010010010000000000010000110001000100011000;
nRam[262] <= 68'b01000000000000000000010000010001100000000000010101000010000010010000;
nRam[263] <= 68'b00100001000000011100010100000000110010000000001110001000100000011000;
nRam[264] <= 68'b00000000000000000000001000000000100000000110000101000000000000000000;
nRam[265] <= 68'b00000110000000000000000000000000000000001000000010000000000000000000;
nRam[266] <= 68'b01000000000000000000010000000000100100001010001100110010000001000000;
nRam[267] <= 68'b01000000000000000000000000000000000100001010001100000000000001000000;
nRam[268] <= 68'b01100001000000011000000000000000100001100010000000000000110000000000;
nRam[269] <= 68'b01000001000000000000010000000000100000000110000101010000000000010000;
nRam[270] <= 68'b00101000000000001000010000001000101010000000000101100000000000100001;
nRam[271] <= 68'b10000110000000000000000000001000001000001000000101100000000000100001;
nRam[272] <= 68'b00000000000000000000000000001000000100000000000001000000000001010001;
nRam[273] <= 68'b00100010000100111000100000000000110010100000000001000000110000010000;
nRam[274] <= 68'b00100100000100111100000000001000000100000000000001000000000001011001;
nRam[275] <= 68'b00100011000000011000010100000000010000000000001110001000100000011000;
nRam[276] <= 68'b00000000000000000000000000011001100110100000010001000000011011010001;
nRam[277] <= 68'b00000000000000000000000000000000000000000000000010000000000000000000;
nRam[278] <= 68'b00000000000100100000010001001000100100000000000001000000011001001001;
nRam[279] <= 68'b00100100001000111100001000000000100010000000000101000000000000010000;
nRam[280] <= 68'b01000001000000000000000000010001100000000010000010000000000000000000;
nRam[281] <= 68'b00100010000000011010000000000000110100000000011110001100100100011000;
nRam[282] <= 68'b11100101000000011100000100000000001000010000010101000000011010000000;
nRam[283] <= 68'b00010000000000000000100000000000100001100010001100000000110000000000;
nRam[284] <= 68'b00100010000100111000010001001000000100000000000000000000000001011001;
nRam[285] <= 68'b00010000000000000010000000000000100100000010001110000000000000011000;
nRam[286] <= 68'b11100011000000011100001000010101100000010000000101000000000000000000;
nRam[287] <= 68'b00100000000000011000000000110010100100011111010001100000000001000000;
nRam[288] <= 68'b10000000000100000000000000001000100110110000000001000000000001011001;
nRam[289] <= 68'b11000001000000000000000000001001000100010000001001000000000011010001;
nRam[290] <= 68'b00100100000100111100000000000000000000000000000101100000000000010000;
nRam[291] <= 68'b10000000000100100000000001001001000100010000001001000000000011001001;
nRam[292] <= 68'b11000001000000000000000000000000000000010000000010000000000000000000;
nRam[293] <= 68'b00110100001100100000000000000000100000000000000101100100000100010000;
nRam[294] <= 68'b00000001000001000000000001000000000000000000000101000000000000010000;
nRam[295] <= 68'b00000001000010000000010001000000100000000000000101000100000010010000;
nRam[296] <= 68'b00100000000100111000000000010000101000010111010101000100000100110010;
nRam[297] <= 68'b11100101000000011100000000000000000000010000000010000000000000000000;
nRam[298] <= 68'b11100101000000011000000000000000100000010000010010000100000100000000;
nRam[299] <= 68'b00000000000000000000000000001000001000000000000101000000000000110001;
nRam[300] <= 68'b00000000000000000000000000000000000000000000000010000000000000000000;
nRam[301] <= 68'b00000000000000000000000000000000000000000000000010000000000000000000;
nRam[302] <= 68'b00000000000000000000000000000000000000000000000010000000000000000000;
nRam[303] <= 68'b00000001000000000000000000001000001001100000000001000000110000110001;
nRam[304] <= 68'b00000001000001000000000001001000000100000000000001010000000001011001;
nRam[305] <= 68'b00100000000000001000001000000000100000000000000010000100000010000000;
nRam[306] <= 68'b11000001000000000000010000001001001000010000000101000000000000110001;
nRam[307] <= 68'b00000000000110000000000001000000100000000000000101000100000100010000;
nRam[308] <= 68'b00000000000101000000000001000000100000000000000101000100000100010000;
nRam[309] <= 68'b00000000000010100000000001010000000100000000000101000000000000010000;
nRam[310] <= 68'b00000000000101000000000001001010000100000000000001010000000001011001;
nRam[311] <= 68'b11100101001000011100000000000000010000010000010010001000000000100000;
nRam[312] <= 68'b00100000000000001000000000001000001000000000000110000000000000110001;
nRam[313] <= 68'b00100000000000011000000000000000100000000100011100000101000100011000;
nRam[314] <= 68'b00100000000000011000000000010000110100000000011100000101000100011000;
nRam[315] <= 68'b01100011100000011000000100010010000000000000000101110000000000000011;
nRam[316] <= 68'b01100010000000011000010100000000010000000000001100000001000000011000;
nRam[317] <= 68'b10000000000100100000000001001000000100010000000001000000000001011001;
nRam[318] <= 68'b01100010000000011000010100000010010000000000001100110001000100011000;
nRam[319] <= 68'b01100011000000011000010000010000000100000000011101110000000001011000;
nRam[320] <= 68'b00000000000000000000010000000000100000000110000101000000000000010000;
nRam[321] <= 68'b00000000000000000000000000000000000000011100001110000000000000011000;
nRam[322] <= 68'b10100000000000001000010000001000101000000110000101000000000000100001;
nRam[323] <= 68'b00100000000000011000000000110001100100001111011001100000000011000010;
nRam[324] <= 68'b00000001000000000000010000000001100001001010000101000010100010010000;
nRam[325] <= 68'b00100010001000111000010000010000000100000000011101000000000001010000;
nRam[326] <= 68'b00100100000100111100000000000000000000000000000101000000000000010000;
nRam[327] <= 68'b00100010000100011000010001010000000100000000011100010000000001010000;
nRam[328] <= 68'b01000001000000000000000100010000011000000000000010000000000000000000;
nRam[329] <= 68'b00000000000000000000010000000000100010000000000101000010001000010000;
nRam[330] <= 68'b00100000000100111000000000000000100000000010000100100000000000010000;
nRam[331] <= 68'b00100010000000011000010000001000001000000000000101000000000000110001;
nRam[332] <= 68'b00000001000000000000010000000000100000000000000101000100000010010000;
nRam[333] <= 68'b00000000000000000000000000000000000000000000000010000000000000000000;
nRam[334] <= 68'b00000000000000000000001000000000100100000000000000110010000001011000;
nRam[335] <= 68'b00000000011000000000000000000010110110000000001100000000001101011000;

	end
	
	always @( posedge clk) nanoOutput <= nRam[ nanoAddr];
endmodule